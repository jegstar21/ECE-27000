(* blackbox *)
module simon #(
  parameter DELAY=2
)(
  input logic clk, reset,
  input logic [19:0] in,
  output logic [7:0] left, right,
  output logic [63:0] ss,
  output logic win, lose
);

// This file is INTENTIONALLY empty!
// Do not enter any code here! - NM

endmodule
